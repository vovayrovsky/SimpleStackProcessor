`timescale 1ns / 1ps

module ALU(
    input wire [2 : 0] func,

    input wire [15 : 0] i0,
    input wire [15 : 0] i1,
    
    output reg [15 : 0] o0
    );


endmodule
